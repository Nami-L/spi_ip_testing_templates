`ifndef SPI_IP_UVC_SEQUENCER_SV
`define SPI_IP_UVC_SEQUENCER_SV


class spi_ip_uvc_sequencer extends uvm_sequencer #(spi_ip_uvc_sequence_item);

  `uvm_component_utils(spi_ip_uvc_sequencer)

  spi_ip_uvc_config m_config;

  extern function new(string name, uvm_component parent);

  extern function void build_phase(uvm_phase phase);

endclass : spi_ip_uvc_sequencer

function spi_ip_uvc_sequencer::new(string name, uvm_component parent);
super.new(name,parent);
endfunction:new

function void spi_ip_uvc_sequencer::build_phase(uvm_phase phase);

if(!uvm_config_db#(spi_ip_uvc_config)::get(get_parent(),"","config",m_config))begin
    `uvm_fatal(get_name(), "Could not retrieve spi_ip_uvc_config from config db")

end
endfunction:build_phase



`endif // SPI_IP_UVC_SEQUENCER_SV
